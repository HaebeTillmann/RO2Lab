`define ALU_ADD 6'b000001
`define ALU_SUB 6'b100001
`define ALU_AND 6'b011101
`define ALU_OR 6'b011001
`define ALU_XOR 6'b010001
`define ALU_SLL 6'b000101
`define ALU_SRA 6'b110101
`define ALU_SRL 6'b00101
`define ALU_SLT 6'b001001
`define ALU_SLTU 6'b001101
`define ALU_EQ 6'b?00010
`define ALU_NE 6'b?00110
`define ALU_LT 6'b?10010
`define ALU_GE 6'b?10110
`define ALU_LTU 6'b?11010
`define ALU_GEU 6'b?11110